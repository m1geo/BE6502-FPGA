module microcode(
    input clk,
    input enable,
    input reset,
    input [8:0] addr,
    output reg [31:0] data );

localparam RESET = 9'b111111111;

reg [31:0] microcode_rom[0:511];

always @(posedge clk)
    if( enable )
        data <= microcode_rom[reset ? RESET : addr];

// Vivado didn't like this. It was unhappy with the $readmemb directive for synthesis. Listing the ROM out worked.
/*initial $readmemb("BE6502-FPGA/be6502_fpga/verilog-65C02-microcode-main/generic/microcode.mem", microcode_rom, 0 );*/

// Not all memory addresses are specified! 
initial begin
    microcode_rom[9'h000] = 32'b10011001011110011001010000011000;
    microcode_rom[9'h001] = 32'b10000011110000000011010000001101;
    microcode_rom[9'h004] = 32'b10000011110000111101010000000010;
    microcode_rom[9'h005] = 32'b10000011110000111011010000000000;
    microcode_rom[9'h006] = 32'b10000011110000111011000000000010;
    microcode_rom[9'h008] = 32'b10011011011110011001010000010110;
    microcode_rom[9'h009] = 32'b10000100010000000000000001001101;
    microcode_rom[9'h00A] = 32'b11000100001100010101000000011011;
    microcode_rom[9'h00C] = 32'b10000100110000111101010000000100;
    microcode_rom[9'h00D] = 32'b10000100110000000011010000000001;
    microcode_rom[9'h00E] = 32'b10000100110000111011000000000100;
    microcode_rom[9'h010] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h011] = 32'b10000011110000111011010000001111;
    microcode_rom[9'h012] = 32'b10000011110000111011010000001101;
    microcode_rom[9'h014] = 32'b10000011110000111110000000000010;
    microcode_rom[9'h015] = 32'b10000011110000000011010000000000;
    microcode_rom[9'h016] = 32'b10000011110000000011000000000010;
    microcode_rom[9'h018] = 32'b10000100000000000000000000000011;
    microcode_rom[9'h019] = 32'b10000100110000000011010000010010;
    microcode_rom[9'h01A] = 32'b11000100001100010001000100011000;
    microcode_rom[9'h01C] = 32'b10000100110000111110000000000100;
    microcode_rom[9'h01D] = 32'b10000100110000000011010000010001;
    microcode_rom[9'h01E] = 32'b10000100110000111011000000000101;
    microcode_rom[9'h020] = 32'b10011001011110011001010000001001;
    microcode_rom[9'h021] = 32'b10000011110000000010110000001101;
    microcode_rom[9'h024] = 32'b10000011110000111010100000000000;
    microcode_rom[9'h025] = 32'b10000011110000111010110000000000;
    microcode_rom[9'h026] = 32'b10000011110000111100100000000010;
    microcode_rom[9'h028] = 32'b10000101011110011001000100010100;
    microcode_rom[9'h029] = 32'b10000100010000000000000001001011;
    microcode_rom[9'h02A] = 32'b11000100001100010101001000011011;
    microcode_rom[9'h02C] = 32'b10000100110000111010100000000001;
    microcode_rom[9'h02D] = 32'b10000100110000000010110000000001;
    microcode_rom[9'h02E] = 32'b10000100110000111100100000000100;
    microcode_rom[9'h030] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h031] = 32'b10000011110000111010110000001111;
    microcode_rom[9'h032] = 32'b10000011110000111010110000001101;
    microcode_rom[9'h034] = 32'b10000011110000000010100000000000;
    microcode_rom[9'h035] = 32'b10000011110000000010110000000000;
    microcode_rom[9'h036] = 32'b10000011110000000100100000000010;
    microcode_rom[9'h038] = 32'b10000100000000111001010100000011;
    microcode_rom[9'h039] = 32'b10000100110000000010110000010010;
    microcode_rom[9'h03A] = 32'b11000100001100010001010000011000;
    microcode_rom[9'h03C] = 32'b10000100110000000010100000010001;
    microcode_rom[9'h03D] = 32'b10000100110000000010110000010001;
    microcode_rom[9'h03E] = 32'b10000100110000111100100000000101;
    microcode_rom[9'h040] = 32'b10000101011110011001000100011100;
    microcode_rom[9'h041] = 32'b10000011110000000010010000001101;
    microcode_rom[9'h045] = 32'b10000011110000111010010000000000;
    microcode_rom[9'h046] = 32'b10000011110000111100110000000010;
    microcode_rom[9'h048] = 32'b10011011011110011001010001000110;
    microcode_rom[9'h049] = 32'b10000100010000000000000001001001;
    microcode_rom[9'h04A] = 32'b11000100001100010111000000011011;
    microcode_rom[9'h04C] = 32'b10000100010000000000000000000110;
    microcode_rom[9'h04D] = 32'b10000100110000000010010000000001;
    microcode_rom[9'h04E] = 32'b10000100110000111100110000000100;
    microcode_rom[9'h050] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h051] = 32'b10000011110000111010010000001111;
    microcode_rom[9'h052] = 32'b10000011110000111010010000001101;
    microcode_rom[9'h055] = 32'b10000011110000000010010000000000;
    microcode_rom[9'h056] = 32'b10000011110000000100110000000010;
    microcode_rom[9'h058] = 32'b10000100000000000000000000100000;
    microcode_rom[9'h059] = 32'b10000100110000000010010000010010;
    microcode_rom[9'h05A] = 32'b10011011011110011001010001001000;
    microcode_rom[9'h05D] = 32'b10000100110000000010010000010001;
    microcode_rom[9'h05E] = 32'b10000100110000111100110000000101;
    microcode_rom[9'h060] = 32'b10000101011110011001000100001011;
    microcode_rom[9'h061] = 32'b10000011110000000000110000001101;
    microcode_rom[9'h064] = 32'b10010011010000111000000001010110;
    microcode_rom[9'h065] = 32'b10000011110000111000110000000000;
    microcode_rom[9'h066] = 32'b10000011110000111101000000000010;
    microcode_rom[9'h068] = 32'b10000101011110011001000100000111;
    microcode_rom[9'h069] = 32'b10000100010000000000000001000011;
    microcode_rom[9'h06A] = 32'b11000100001100010111001000011011;
    microcode_rom[9'h06C] = 32'b10000100010000000000110000100111;
    microcode_rom[9'h07C] = 32'b10000100010000000000110000101101;
    microcode_rom[9'h06D] = 32'b10000100110000000000110000000001;
    microcode_rom[9'h06E] = 32'b10000100110000111101000000000100;
    microcode_rom[9'h070] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h071] = 32'b10000011110000111000110000001111;
    microcode_rom[9'h072] = 32'b10000011110000111000110000001101;
    microcode_rom[9'h074] = 32'b10010011010000000000000001010110;
    microcode_rom[9'h075] = 32'b10000011110000000000110000000000;
    microcode_rom[9'h076] = 32'b10000011110000000101000000000010;
    microcode_rom[9'h078] = 32'b10000100000000000000000000100000;
    microcode_rom[9'h079] = 32'b10000100110000000000110000010010;
    microcode_rom[9'h07A] = 32'b10000101011110011001000100010011;
    microcode_rom[9'h07D] = 32'b10000100110000000000110000010001;
    microcode_rom[9'h07E] = 32'b10000100110000111101000000000101;
    microcode_rom[9'h080] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h081] = 32'b10000011110000000001100000100011;
    microcode_rom[9'h084] = 32'b10010011010000111000000001001000;
    microcode_rom[9'h085] = 32'b10010011010000111000000001000110;
    microcode_rom[9'h086] = 32'b10010011010000111000000001000111;
    microcode_rom[9'h088] = 32'b11000100001010001001010000011000;
    microcode_rom[9'h089] = 32'b10000100010000000000000001010111;
    microcode_rom[9'h08A] = 32'b11000100001100000001000000011000;
    microcode_rom[9'h08C] = 32'b10000100110000111010000000100000;
    microcode_rom[9'h08D] = 32'b10000100110000111001100000100000;
    microcode_rom[9'h08E] = 32'b10000100110000111001110000100000;
    microcode_rom[9'h090] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h091] = 32'b10000011110000111001100000100101;
    microcode_rom[9'h092] = 32'b10000011110000111001100000100011;
    microcode_rom[9'h094] = 32'b10010011010000000000000001001000;
    microcode_rom[9'h095] = 32'b10010011010000000000000001000110;
    microcode_rom[9'h096] = 32'b10010011010000001000000001000111;
    microcode_rom[9'h098] = 32'b11000100001100001001000000011000;
    microcode_rom[9'h099] = 32'b10000100110000111001100000100010;
    microcode_rom[9'h09A] = 32'b10000100001110000001000000000000;
    microcode_rom[9'h09C] = 32'b10000100110000111101100000100000;
    microcode_rom[9'h09D] = 32'b10000100110000111001100000100001;
    microcode_rom[9'h09E] = 32'b10000100110000111101100000100001;
    microcode_rom[9'h0A0] = 32'b10000100010000000000000001000010;
    microcode_rom[9'h0A1] = 32'b10000011110000000000000000001101;
    microcode_rom[9'h0A2] = 32'b10000100010000000000000001000001;
    microcode_rom[9'h0A4] = 32'b10000011110000111000100000000000;
    microcode_rom[9'h0A5] = 32'b10000011110000111000000000000000;
    microcode_rom[9'h0A6] = 32'b10000011110000111000010000000000;
    microcode_rom[9'h0A8] = 32'b11000100001010010001000000011000;
    microcode_rom[9'h0A9] = 32'b10000100010000000000000001000000;
    microcode_rom[9'h0AA] = 32'b11000100001000010001000000011000;
    microcode_rom[9'h0AC] = 32'b10000100110000000000100000000001;
    microcode_rom[9'h0AD] = 32'b10000100110000000000000000000001;
    microcode_rom[9'h0AE] = 32'b10000100110000000000010000000001;
    microcode_rom[9'h0B0] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h0B1] = 32'b10000011110000111000000000001111;
    microcode_rom[9'h0B2] = 32'b10000011110000111000000000001101;
    microcode_rom[9'h0B4] = 32'b10000011110000000000100000000000;
    microcode_rom[9'h0B5] = 32'b10000011110000000000000000000000;
    microcode_rom[9'h0B6] = 32'b10000011110000001000010000000000;
    microcode_rom[9'h0B8] = 32'b10000100000000111000110010000000;
    microcode_rom[9'h0B9] = 32'b10000100110000000000000000010010;
    microcode_rom[9'h0BA] = 32'b11000100001000011001000000011000;
    microcode_rom[9'h0BC] = 32'b10000100110000000000100000010001;
    microcode_rom[9'h0BD] = 32'b10000100110000000000000000010001;
    microcode_rom[9'h0BE] = 32'b10000100110000000000010000010010;
    microcode_rom[9'h0C0] = 32'b10000100010000000000000001010001;
    microcode_rom[9'h0C1] = 32'b10000011110000000011100000001101;
    microcode_rom[9'h0C4] = 32'b10000011110000111100010000000000;
    microcode_rom[9'h0C5] = 32'b10000011110000111011100000000000;
    microcode_rom[9'h0C6] = 32'b10000011110000111001010000000010;
    microcode_rom[9'h0C8] = 32'b11000100001010001001000100011000;
    microcode_rom[9'h0C9] = 32'b10000100010000000000000001001110;
    microcode_rom[9'h0CA] = 32'b11000100001000000001010000011000;
    microcode_rom[9'h0CC] = 32'b10000100110000111100010000000001;
    microcode_rom[9'h0CD] = 32'b10000100110000000011100000000001;
    microcode_rom[9'h0CE] = 32'b10000100110000111001010000000100;
    microcode_rom[9'h0D0] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h0D1] = 32'b10000011110000111011100000001111;
    microcode_rom[9'h0D2] = 32'b10000011110000111011100000001101;
    microcode_rom[9'h0D5] = 32'b10000011110000000011100000000000;
    microcode_rom[9'h0D6] = 32'b10000011110000000001010000000010;
    microcode_rom[9'h0D8] = 32'b10000100000000000000000001000000;
    microcode_rom[9'h0D9] = 32'b10000100110000000011100000010010;
    microcode_rom[9'h0DA] = 32'b10011011011110011001010001000111;
    microcode_rom[9'h0DD] = 32'b10000100110000000011100000010001;
    microcode_rom[9'h0DE] = 32'b10000100110000111001010000000101;
    microcode_rom[9'h0E0] = 32'b10000100010000000000000001010000;
    microcode_rom[9'h0E1] = 32'b10000011110000000011110000001101;
    microcode_rom[9'h0E4] = 32'b10000011110000111100000000000000;
    microcode_rom[9'h0E5] = 32'b10000011110000111011110000000000;
    microcode_rom[9'h0E6] = 32'b10000011110000111001000000000010;
    microcode_rom[9'h0E8] = 32'b11000100001000000001000100011000;
    microcode_rom[9'h0E9] = 32'b10000100010000000000000001001111;
    microcode_rom[9'h0EA] = 32'b10000100000000000000000000000000;
    microcode_rom[9'h0EC] = 32'b10000100110000111100000000000001;
    microcode_rom[9'h0ED] = 32'b10000100110000000011110000000001;
    microcode_rom[9'h0EE] = 32'b10000100110000111001000000000100;
    microcode_rom[9'h0F0] = 32'b10000111010000000000000000000011;
    microcode_rom[9'h0F1] = 32'b10000011110000111011110000001111;
    microcode_rom[9'h0F2] = 32'b10000011110000111011110000001101;
    microcode_rom[9'h0F5] = 32'b10000011110000000011110000000000;
    microcode_rom[9'h0F6] = 32'b10000011110000000001000000000010;
    microcode_rom[9'h0F8] = 32'b10000100000000000000000001000000;
    microcode_rom[9'h0F9] = 32'b10000100110000000011110000010010;
    microcode_rom[9'h0FA] = 32'b10000101011110011001000100001000;
    microcode_rom[9'h0FD] = 32'b10000100110000000011110000010001;
    microcode_rom[9'h0FE] = 32'b10000100110000111001000000000101;
    microcode_rom[9'h100] = 32'b10000001100000000000000000000000;
    microcode_rom[9'h101] = 32'b10000010010000111000000000000000;
    microcode_rom[9'h102] = 32'b10010000100000000000000000000000;
    microcode_rom[9'h103] = 32'b10000100000000000000000000000000;
    microcode_rom[9'h104] = 32'b10000010010000111000000000000010;
    microcode_rom[9'h105] = 32'b10000010010000000000000000000010;
    microcode_rom[9'h106] = 32'b10000010010000111000000000000011;
    microcode_rom[9'h107] = 32'b10000001010000000000000001000000;
    microcode_rom[9'h108] = 32'b10000001010000000000000001000001;
    microcode_rom[9'h109] = 32'b11111000011110011001010000001010;
    microcode_rom[9'h10A] = 32'b11000001010000000000000000000110;
    microcode_rom[9'h10B] = 32'b10000101011110011001000100001100;
    microcode_rom[9'h10C] = 32'b10001110010000111000000000000011;
    microcode_rom[9'h10D] = 32'b10001100010000000000000000001110;
    microcode_rom[9'h10E] = 32'b10001010010000111000000000000000;
    microcode_rom[9'h10F] = 32'b10001100010000000000000000010000;
    microcode_rom[9'h110] = 32'b10001010010000001000000000000000;
    microcode_rom[9'h111] = 32'b10000010010000000000000000000000;
    microcode_rom[9'h112] = 32'b10000010010000001000000000000000;
    microcode_rom[9'h113] = 32'b10000001010000000000000001000010;
    microcode_rom[9'h114] = 32'b10000001010000000000000000010101;
    microcode_rom[9'h115] = 32'b10100100000000111110110010010111;
    microcode_rom[9'h116] = 32'b10100001010000000000000100000011;
    microcode_rom[9'h117] = 32'b11000100000000111000110100011000;
    microcode_rom[9'h118] = 32'b11111000011110011001010000011001;
    microcode_rom[9'h119] = 32'b11011000011110011001010000011010;
    microcode_rom[9'h11A] = 32'b10101111010001010000000100011011;
    microcode_rom[9'h11B] = 32'b10001100010000000000000000101000;
    microcode_rom[9'h11C] = 32'b10000101011110011001000100011101;
    microcode_rom[9'h11D] = 32'b00000101011110011001000100011110;
    microcode_rom[9'h11E] = 32'b00000010010000111110110000010101;
    microcode_rom[9'h120] = 32'b10010010100000111000000000000000;
    microcode_rom[9'h121] = 32'b10010010100000000000000000000000;
    microcode_rom[9'h122] = 32'b10010010100000001000000000000000;
    microcode_rom[9'h123] = 32'b10001100010000000000000000100100;
    microcode_rom[9'h124] = 32'b10011010100000111000000000000000;
    microcode_rom[9'h125] = 32'b10001100010000000000000000100110;
    microcode_rom[9'h126] = 32'b10011010100000001000000000000000;
    microcode_rom[9'h127] = 32'b10000010010000111000000000101110;
    microcode_rom[9'h128] = 32'b10000010010000111000000000101001;
    microcode_rom[9'h129] = 32'b10000100000000000000000001100000;
    microcode_rom[9'h12A] = 32'b11000100000000010000010000000000;
    microcode_rom[9'h12B] = 32'b11000100000000110000110000011000;
    microcode_rom[9'h12C] = 32'b11000100000000111100110000011011;
    microcode_rom[9'h12D] = 32'b10000010010000000000000000101110;
    microcode_rom[9'h12E] = 32'b10001100010000000000000000101111;
    microcode_rom[9'h12F] = 32'b10000010010000111000000000110000;
    microcode_rom[9'h130] = 32'b10000100000000000000000000000000;
    microcode_rom[9'h131] = 32'b11000100000000111100111000011011;
    microcode_rom[9'h132] = 32'b11000100000000111110110000011011;
    microcode_rom[9'h133] = 32'b11000100000000111110111000011011;
    microcode_rom[9'h140] = 32'b11000100001100111000000000011000;
    microcode_rom[9'h141] = 32'b11000100001000111000000000011000;
    microcode_rom[9'h142] = 32'b11000100001010111000000000011000;
    microcode_rom[9'h143] = 32'b11000100001100010000111110011011;
    microcode_rom[9'h144] = 32'b00000001010000111000110100010111;
    microcode_rom[9'h145] = 32'b00000001010000110000110000101011;
    microcode_rom[9'h146] = 32'b10000001010000010001000000000011;
    microcode_rom[9'h147] = 32'b10000001010000000001000000000011;
    microcode_rom[9'h148] = 32'b10000001010000001001000000000011;
    microcode_rom[9'h149] = 32'b11000100001100010000100000011000;
    microcode_rom[9'h14A] = 32'b11100100000000010000010010001000;
    microcode_rom[9'h14B] = 32'b11000100001100010000010000011000;
    microcode_rom[9'h14C] = 32'b00000001010000111100110000101100;
    microcode_rom[9'h14D] = 32'b11000100001100010000000000011000;
    microcode_rom[9'h14E] = 32'b11000100000000010001100100011011;
    microcode_rom[9'h14F] = 32'b11000100001100010001101110011011;
    microcode_rom[9'h150] = 32'b11000100000000000001100100011011;
    microcode_rom[9'h151] = 32'b11000100000000001001100100011011;
    microcode_rom[9'h152] = 32'b00000001010000111100111000110001;
    microcode_rom[9'h153] = 32'b00000001010000111110110000110010;
    microcode_rom[9'h154] = 32'b00000001010000111110111000110011;
    microcode_rom[9'h155] = 32'b00000001010000010000000000101010;
    microcode_rom[9'h156] = 32'b10000001010000111001000000000011;
    microcode_rom[9'h157] = 32'b11100100000000010000010000000000;
    microcode_rom[9'h158] = 32'b00000001010000010001110000101010;
    microcode_rom[9'h160] = 32'b10011000011110011001010001100001;
    microcode_rom[9'h161] = 32'b11111000011110011001010001100010;
    microcode_rom[9'h162] = 32'b11011000011110011001010001100011;
    microcode_rom[9'h163] = 32'b10101111010001010000000001100100;
    microcode_rom[9'h164] = 32'b10001100010000000000000001100101;
    microcode_rom[9'h165] = 32'b10001010010000111000000001100110;
    microcode_rom[9'h166] = 32'b10000100000000111000000001100000;
    microcode_rom[9'h168] = 32'b11111000011110011001010001101001;
    microcode_rom[9'h169] = 32'b11011000011110011001010001101010;
    microcode_rom[9'h16A] = 32'b10101111010001000000000001101011;
    microcode_rom[9'h16B] = 32'b10001100010000000000000001101100;
    microcode_rom[9'h16C] = 32'b10001010010000111000000001101101;
    microcode_rom[9'h16D] = 32'b10000100000000111000000001100000;
    microcode_rom[9'h170] = 32'b10001111010001001000000001110001;
    microcode_rom[9'h171] = 32'b10000100010000111000000001110010;
    microcode_rom[9'h172] = 32'b10000010010000111000000001110011;
    microcode_rom[9'h173] = 32'b10000100000000111000000001110000;
    microcode_rom[9'h180] = 32'b10000001100000000000000000000000;
    microcode_rom[9'h181] = 32'b10000010010000111000000000000000;
    microcode_rom[9'h182] = 32'b10010000100000000000000000000000;
    microcode_rom[9'h183] = 32'b10000100000000000000000000000000;
    microcode_rom[9'h184] = 32'b10000010010000111000000000000010;
    microcode_rom[9'h185] = 32'b10000010010000000000000000000010;
    microcode_rom[9'h186] = 32'b10000010010000111000000000000011;
    microcode_rom[9'h187] = 32'b10000001010000000000000001000000;
    microcode_rom[9'h188] = 32'b10000001010000000000000001000001;
    microcode_rom[9'h189] = 32'b11111000011110011001010000001010;
    microcode_rom[9'h18A] = 32'b11000001010000000000000000000110;
    microcode_rom[9'h18B] = 32'b10000101011110011001000100001100;
    microcode_rom[9'h18C] = 32'b10001110010000111000000000000011;
    microcode_rom[9'h18D] = 32'b10001100010000000000000000001110;
    microcode_rom[9'h18E] = 32'b10001010010000111000000000000000;
    microcode_rom[9'h18F] = 32'b10001100010000000000000000010000;
    microcode_rom[9'h190] = 32'b10001010010000001000000000000000;
    microcode_rom[9'h191] = 32'b10000010010000000000000000000000;
    microcode_rom[9'h192] = 32'b10000010010000001000000000000000;
    microcode_rom[9'h193] = 32'b10000001010000000000000001000010;
    microcode_rom[9'h194] = 32'b10000001010000000000000000010101;
    microcode_rom[9'h195] = 32'b10100100000000111110110010010111;
    microcode_rom[9'h196] = 32'b10100001010000000000000100000011;
    microcode_rom[9'h197] = 32'b11000100000000111000110100011000;
    microcode_rom[9'h198] = 32'b11111000011110011001010000011001;
    microcode_rom[9'h199] = 32'b11011000011110011001010000011010;
    microcode_rom[9'h19A] = 32'b10101111010001010000000100011011;
    microcode_rom[9'h19B] = 32'b10001100010000000000000000101000;
    microcode_rom[9'h19C] = 32'b10000101011110011001000100011101;
    microcode_rom[9'h19D] = 32'b00000101011110011001000100011110;
    microcode_rom[9'h19E] = 32'b00000010010000111110110000010101;
    microcode_rom[9'h1A0] = 32'b10010010100000111000000000000000;
    microcode_rom[9'h1A1] = 32'b10010010100000000000000000000000;
    microcode_rom[9'h1A2] = 32'b10010010100000001000000000000000;
    microcode_rom[9'h1A3] = 32'b10001100010000000000000000100100;
    microcode_rom[9'h1A4] = 32'b10011010100000111000000000000000;
    microcode_rom[9'h1A5] = 32'b10001100010000000000000000100110;
    microcode_rom[9'h1A6] = 32'b10011010100000001000000000000000;
    microcode_rom[9'h1A7] = 32'b10000010010000111000000000101110;
    microcode_rom[9'h1A8] = 32'b10000010010000111000000000101001;
    microcode_rom[9'h1A9] = 32'b10000100000000000000000001100000;
    microcode_rom[9'h1AA] = 32'b11000100000000010000010000000000;
    microcode_rom[9'h1AB] = 32'b11000100000000110000110000011000;
    microcode_rom[9'h1AC] = 32'b11000100000000111100110000011011;
    microcode_rom[9'h1AD] = 32'b10000010010000000000000000101110;
    microcode_rom[9'h1AE] = 32'b10001100010000000000000000101111;
    microcode_rom[9'h1AF] = 32'b10000010010000111000000000110000;
    microcode_rom[9'h1B0] = 32'b10000100000000000000000000000000;
    microcode_rom[9'h1B1] = 32'b11000100000000111100111000011011;
    microcode_rom[9'h1B2] = 32'b11000100000000111110110000011011;
    microcode_rom[9'h1B3] = 32'b11000100000000111110111000011011;
    microcode_rom[9'h1C0] = 32'b11000100001100111000000000011000;
    microcode_rom[9'h1C1] = 32'b11000100001000111000000000011000;
    microcode_rom[9'h1C2] = 32'b11000100001010111000000000011000;
    microcode_rom[9'h1C3] = 32'b11000000011100010000111111011001;
    microcode_rom[9'h1C4] = 32'b00000001010000111000110100010111;
    microcode_rom[9'h1C5] = 32'b00000001010000110000110000101011;
    microcode_rom[9'h1C6] = 32'b10000001010000010001000000000011;
    microcode_rom[9'h1C7] = 32'b10000001010000000001000000000011;
    microcode_rom[9'h1C8] = 32'b10000001010000001001000000000011;
    microcode_rom[9'h1C9] = 32'b11000100001100010000100000011000;
    microcode_rom[9'h1CA] = 32'b11100100000000010000010010001000;
    microcode_rom[9'h1CB] = 32'b11000100001100010000010000011000;
    microcode_rom[9'h1CC] = 32'b00000001010000111100110000101100;
    microcode_rom[9'h1CD] = 32'b11000100001100010000000000011000;
    microcode_rom[9'h1CE] = 32'b11000100000000010001100100011011;
    microcode_rom[9'h1CF] = 32'b11000000011100010001101111011010;
    microcode_rom[9'h1D0] = 32'b11000100000000000001100100011011;
    microcode_rom[9'h1D1] = 32'b11000100000000001001100100011011;
    microcode_rom[9'h1D2] = 32'b00000001010000111100111000110001;
    microcode_rom[9'h1D3] = 32'b00000001010000111110110000110010;
    microcode_rom[9'h1D4] = 32'b00000001010000111110111000110011;
    microcode_rom[9'h1D5] = 32'b00000001010000010000000000101010;
    microcode_rom[9'h1D6] = 32'b10000001010000111001000000000011;
    microcode_rom[9'h1D7] = 32'b11100100000000010000010000000000;
    microcode_rom[9'h1D8] = 32'b00000001010000010001110000101010;
    microcode_rom[9'h1D9] = 32'b11000100001100010000110000011011;
    microcode_rom[9'h1DA] = 32'b11000100001100010001100100011011;
    microcode_rom[9'h1E0] = 32'b10011000011110011001010001101000;
    microcode_rom[9'h1E1] = 32'b11111000011110011001010001100010;
    microcode_rom[9'h1E2] = 32'b11011000011110011001010001100011;
    microcode_rom[9'h1E3] = 32'b10101111010001010000000001100100;
    microcode_rom[9'h1E4] = 32'b10001100010000000000000001100101;
    microcode_rom[9'h1E5] = 32'b10001010010000111000000001100110;
    microcode_rom[9'h1E6] = 32'b10000100000000111000000001100000;
    microcode_rom[9'h1E8] = 32'b11111000011110011001010001101001;
    microcode_rom[9'h1E9] = 32'b11011000011110011001010001101010;
    microcode_rom[9'h1EA] = 32'b10101111010001000000000001101011;
    microcode_rom[9'h1EB] = 32'b10001100010000000000000001101100;
    microcode_rom[9'h1EC] = 32'b10001010010000111000000001101101;
    microcode_rom[9'h1ED] = 32'b10000100000000111000000001100000;
    microcode_rom[9'h1F0] = 32'b10001111010001001000000001110001;
    microcode_rom[9'h1F1] = 32'b10000100010000111000000001110010;
    microcode_rom[9'h1F2] = 32'b10000010010000111000000001110011;
    microcode_rom[9'h1F3] = 32'b10000100000000111000000001110000;
    microcode_rom[9'h1FF] = 32'b00000000010000000000000001110000;
end

endmodule